magic
tech sky130A
magscale 1 2
timestamp 1768503958
<< error_s >>
rect 288 -190 294 -9
rect 288 -196 447 -190
<< locali >>
rect 152 1968 859 2040
rect -200 -9 1400 0
rect -200 -196 288 -9
rect 447 -196 1400 -9
rect -200 -200 1400 -196
<< viali >>
rect 288 -196 447 -9
<< metal1 >>
rect 160 39 224 3960
rect 672 3761 1166 3953
rect 288 680 459 3312
rect 974 3050 1166 3761
rect 683 2858 1166 3050
rect 974 1433 1166 2858
rect 707 1241 1166 1433
rect 288 600 480 680
rect 288 -9 459 600
rect 974 507 1166 1241
rect 695 315 1166 507
rect 672 40 864 120
rect 447 -196 459 -9
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1768503958
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1> ../JNW_ATR_SKY130A
timestamp 1768503958
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1 ../JNW_ATR_SKY130A
timestamp 1768503958
transform 1 0 0 0 1 1600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<0> ../JNW_ATR_SKY130A
timestamp 1768503958
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<1> ../JNW_ATR_SKY130A
timestamp 1768503958
transform 1 0 0 0 1 3200
box -184 -128 1336 928
<< labels >>
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 1 nsew signal bidirectional
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
